** sch_path: /foss/designs/asitic-example/examples/sq_1nH_2.5GHz/xschem/tb-ind.sch
**.subckt tb-ind
V1 p1 GND DC 0 AC 1
x1 p1 GND GND l0
**** begin user architecture code

.ac lin 100k 100Meg 40G
.control
destroy all
run
save all
let z_complex = -v(p1)/i(v1)
let z = mag(z_complex)
let x = imag(z_complex)
let r = real(z_complex)
write tb-impedance.raw
plot z x r
.endc

.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt
**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/asitic-example/examples/sq_1nH_2.5GHz/xschem/l0.sym # of pins=3
** sym_path: /foss/designs/asitic-example/examples/sq_1nH_2.5GHz/xschem/l0.sym
** sch_path: /foss/designs/asitic-example/examples/sq_1nH_2.5GHz/xschem/l0.sch
.subckt l0 p1 p2 sub
*.iopin sub
*.iopin p1
*.iopin p2
R net2 p2 2.857 m=1
L p1 net2 1.006n m=1
Rs1 net1 sub 27.37 m=1
Cs1 p1 net1 33.97f m=1
Cs2 p2 net3 36.78f m=1
Rs2 net3 sub -9 m=1
.ends

.GLOBAL GND
.end
