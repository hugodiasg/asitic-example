magic
tech sky130A
magscale 1 2
timestamp 1726236408
<< metal4 >>
rect -5358 4699 -200 4740
rect -5358 161 -456 4699
rect -220 161 -200 4699
rect -5358 120 -200 161
rect 200 4699 5358 4740
rect 200 161 5102 4699
rect 5338 161 5358 4699
rect 200 120 5358 161
rect -5358 -161 -200 -120
rect -5358 -4699 -456 -161
rect -220 -4699 -200 -161
rect -5358 -4740 -200 -4699
rect 200 -161 5358 -120
rect 200 -4699 5102 -161
rect 5338 -4699 5358 -161
rect 200 -4740 5358 -4699
<< via4 >>
rect -456 161 -220 4699
rect 5102 161 5338 4699
rect -456 -4699 -220 -161
rect 5102 -4699 5338 -161
<< mimcap2 >>
rect -5278 4620 -818 4660
rect -5278 240 -5238 4620
rect -858 240 -818 4620
rect -5278 200 -818 240
rect 280 4620 4740 4660
rect 280 240 320 4620
rect 4700 240 4740 4620
rect 280 200 4740 240
rect -5278 -240 -818 -200
rect -5278 -4620 -5238 -240
rect -858 -4620 -818 -240
rect -5278 -4660 -818 -4620
rect 280 -240 4740 -200
rect 280 -4620 320 -240
rect 4700 -4620 4740 -240
rect 280 -4660 4740 -4620
<< mimcap2contact >>
rect -5238 240 -858 4620
rect 320 240 4700 4620
rect -5238 -4620 -858 -240
rect 320 -4620 4700 -240
<< metal5 >>
rect -3208 4644 -2888 4860
rect -498 4699 -178 4860
rect -5262 4620 -834 4644
rect -5262 240 -5238 4620
rect -858 240 -834 4620
rect -5262 216 -834 240
rect -3208 -216 -2888 216
rect -498 161 -456 4699
rect -220 161 -178 4699
rect 2350 4644 2670 4860
rect 5060 4699 5380 4860
rect 296 4620 4724 4644
rect 296 240 320 4620
rect 4700 240 4724 4620
rect 296 216 4724 240
rect -498 -161 -178 161
rect -5262 -240 -834 -216
rect -5262 -4620 -5238 -240
rect -858 -4620 -834 -240
rect -5262 -4644 -834 -4620
rect -3208 -4860 -2888 -4644
rect -498 -4699 -456 -161
rect -220 -4699 -178 -161
rect 2350 -216 2670 216
rect 5060 161 5102 4699
rect 5338 161 5380 4699
rect 5060 -161 5380 161
rect 296 -240 4724 -216
rect 296 -4620 320 -240
rect 4700 -4620 4724 -240
rect 296 -4644 4724 -4620
rect -498 -4860 -178 -4699
rect 2350 -4860 2670 -4644
rect 5060 -4699 5102 -161
rect 5338 -4699 5380 -161
rect 5060 -4860 5380 -4699
<< properties >>
string FIXED_BBOX 200 120 4820 4740
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 22.3 l 22.3 val 1.011k carea 2.00 cperi 0.19 nx 2 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
