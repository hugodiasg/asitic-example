** sch_path: /foss/designs/asitic-example/examples/sq_1nH_2.5GHz/xschem/tb-tran.sch
**.subckt tb-tran
V1 net1 GND sin(0 1.8 2.5G)
V2 v1 net1 0
x1 v1 GND net2 l0
**** begin user architecture code

.tran 0.4p 400p
.control
destroy all
run
let i1 = -i(v2)
plot v1 i1

.endc

.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt
**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/asitic-example/examples/sq_1nH_2.5GHz/xschem/l0.sym # of pins=3
** sym_path: /foss/designs/asitic-example/examples/sq_1nH_2.5GHz/xschem/l0.sym
** sch_path: /foss/designs/asitic-example/examples/sq_1nH_2.5GHz/xschem/l0.sch
.subckt l0 p1 p2 sub
*.iopin sub
*.iopin p1
*.iopin p2
R net2 p2 2.857 m=1
L p1 net2 1.006n m=1
Rs1 net1 sub 27.37 m=1
Cs1 p1 net1 33.97f m=1
Cs2 p2 net3 36.78f m=1
Rs2 net3 sub -9 m=1
.ends

.GLOBAL GND
.end
