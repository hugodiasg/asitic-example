magic
tech sky130A
timestamp 1725456507
<< metal4 >>
rect 26200 24938 27400 25000
rect 26200 23860 26260 24938
rect 27338 23860 27400 24938
rect 26200 18400 27400 23860
<< via4 >>
rect 26260 23860 27338 24938
<< metal5 >>
rect 19600 30400 31600 31600
rect 19600 29000 30200 30200
rect 19600 20800 20800 29000
rect 21000 27600 28800 28800
rect 21000 22200 22200 27600
rect 22400 26200 27400 27400
rect 22400 23600 23600 26200
rect 26200 24938 27400 26200
rect 26200 23860 26260 24938
rect 27338 23860 27400 24938
rect 26200 23800 27400 23860
rect 27600 23600 28800 27600
rect 22400 22400 28800 23600
rect 29000 22200 30200 29000
rect 21000 21000 30200 22200
rect 30400 20800 31600 30400
rect 19600 19600 31600 20800
<< end >>
