magic
tech sky130A
magscale 1 2
timestamp 1726351381
<< psubdiff >>
rect 22876 36800 22900 38800
rect 25200 36800 25224 38800
<< psubdiffcont >>
rect 22900 36800 25200 38800
<< locali >>
rect 25200 36800 25216 38800
<< viali >>
rect 22600 38800 25200 38900
rect 22600 36800 22900 38800
rect 22900 36800 25200 38800
rect 22600 36500 25200 36800
<< metal1 >>
rect 22588 38900 25212 38906
rect 22588 36500 22600 38900
rect 25200 36500 25212 38900
rect 22588 36494 25212 36500
<< via1 >>
rect 22600 36500 25200 38900
<< metal2 >>
rect 22600 38900 25200 38910
rect 22600 36490 25200 36500
<< via2 >>
rect 22600 36500 25200 38900
<< metal3 >>
rect 22590 38900 25210 38905
rect 22590 36500 22600 38900
rect 25200 36500 25210 38900
rect 22590 36495 25210 36500
rect 22800 33600 25200 36495
<< metal4 >>
rect 25400 52450 26500 55100
rect 30950 52450 32050 55150
rect 25400 51350 32050 52450
rect 29000 38900 31400 51350
rect 52200 38900 54600 43400
rect 29000 36500 54600 38900
rect 39200 33600 41600 36500
<< metal5 >>
rect 34700 67400 37100 70300
rect 31000 66900 38000 67400
rect 25600 65900 38000 66900
rect 25600 63000 26600 65900
rect 30900 65000 38000 65900
rect 38200 65000 41500 67400
rect 30900 63300 31900 65000
<< rm5 >>
rect 38000 65000 38200 67400
use l0  l0_0
timestamp 1726236534
transform 1 0 -200 0 1 4200
box 39200 36800 63200 63200
use sky130_fd_pr__cap_mim_m3_2_5YW5FM  sky130_fd_pr__cap_mim_m3_2_5YW5FM_0
timestamp 1726236408
transform 1 0 28958 0 1 59260
box -5358 -4860 5380 4860
<< labels >>
flabel metal5 35400 68700 36500 69800 0 FreeSans 16000 0 0 0 p1
port 1 nsew
flabel metal4 39400 34500 40900 35100 0 FreeSans 16000 0 0 0 p2
port 3 nsew
flabel metal3 23300 34100 24500 35700 0 FreeSans 16000 0 0 0 gnd
port 6 nsew
<< end >>
